library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Logic is port (
	
	hex_A : in std_logic_vector(3 downto 0);
	hex_B : in std_logic_vector(3 downto 0);
	LOG3res : out std_logic_vector(3 downto 0);
);
end Adder;

architecture Behavioural of Logic is 

begin 

with 


end architecture Logic; 